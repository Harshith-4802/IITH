Full wave 5V

V1 0 1 sin(0 5 100 0 0)
D1 1 2 diode
D2 0 2 diode
D3 3 0 diode
D4 3 1 diode
.model diode d(VJ=0.65)
R1 2 3 1k

.control
set color0 = white
set color1 = black

tran 1m 20m 0
plot v(1),v(2,3)
.endc