XOR with NOR GATEs

.subckt nor 1 2 3 4
*1 = Vin1
*2 = Vin2
*3 = Output
*4 = Vdd
m1 5 1 4 4 p1
m2 3 2 5 4 p1
.model p1 PMOS W=10u
m3 3 2 0 0 n1
m4 3 1 0 0 n1
.model n1 NMOS W=1u
.ends nor

Vdd 8 0 dc 5v
Vin1 1 0 DC 5 PULSE(5 0 0 5ns 5ns 100ns 200ns)
Vin2 2 0 DC 5 PULSE(5 0 0 5ns 5ns 50ns 150ns)
X1 1 1 3 8 nor
X2 2 2 4 8 nor
X3 1 2 6 8 nor
X4 3 4 5 8 nor
X5 5 6 7 8 nor

.control
set color0 = white
tran 0.1n 0.2u 0
plot V(1), 6 + V(2), 12 + V(7),18 + V(5)
set xbrushwidth = 2
.endc
