OR GATE

.subckt nor 1 2 3 4
*1 = Vin1
*2 = Vin2
*3 = Output
*4 = Vdd
m1 5 1 4 4 p1
m2 3 2 5 4 p1
.model p1 PMOS W=10u
m3 3 2 0 0 n1
m4 3 1 0 0 n1
.model n1 NMOS W=1u
.ends nor


.subckt not 1 2 3
*1 = Vin
*2 = Vo
*3 = Vdd
m1 2 1 3 3 p1
.model p1 PMOS W=10u
m2 2 1 0 0 n1
.model n1 NMOS W=1u
.ends not


Vdd 4 0 dc 5v
Vin1 1 0 DC 5 PULSE(0 5 0 0.1ns 0.1ns 50ns 100ns)
Vin2 2 0 DC 5 PULSE(0 5 0 0.1ns 0.1ns 100ns 200ns)
X1 1 2 3 4 nor
X2 3 5 4 not

.control
set color0 = white
tran 0.1n 0.2u 0
plot V(1), 6 + V(2), 12 + V(5)
set xbrushwidth = 2
.endc
