NOT GATE

*1 = Vin
*2 = Vo
*3 = Vdd

Vin 1 0 0
m1 2 1 3 3 p1
.model p1 PMOS W=10u
m2 2 1 0 0 n1
.model n1 NMOS W=1u
Vdd 3 0 dc 5v

.control
dc Vin 0 5 0.01
set color0 = white
plot v(2)
set xbrushwidth = 2
.endc
